module cod ( 
	i,
	c
	) ;

input [7:0] i;
inout [2:0] c;
