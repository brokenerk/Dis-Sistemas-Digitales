module sec ( 
	clr,
	clk,
	ent,
	display
	) ;

input  clr;
input  clk;
input [5:0] ent;
inout [6:0] display;
