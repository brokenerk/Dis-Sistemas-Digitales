module ffd ( 
	pre,
	clr,
	clk,
	d,
	q,
	nq
	) ;

input  pre;
input  clr;
input  clk;
input  d;
inout  q;
inout  nq;
