module displays ( 
	r,
	dr
	) ;

input [1:0] r;
inout [6:0] dr;
