LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CONDEC IS
	PORT(CLK, CLR : IN STD_LOGIC;
			C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			E: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			DISPLAY: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);

ATTRIBUTE PIN_NUMBERS OF CONDEC : ENTITY IS
"CLK:1 CLR:2 C(1):3 C(0):4 E(3):5 E(2):6 E(1):7 E(0):8";
END ENTITY;
ARCHITECTURE A_CONDEC OF CONDEC IS
	CONSTANT DIG0 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1000000";
	CONSTANT DIG1 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1111001";
	CONSTANT DIG2 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100100";  
	CONSTANT DIG3 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0110000";
	CONSTANT DIG4 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0011001";
	CONSTANT DIG5 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0010010";
	CONSTANT DIG6 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000010";
	CONSTANT DIG7 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1111000";
	CONSTANT DIG8 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000000";
	CONSTANT DIG9 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0010000";
	CONSTANT APAG : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1111111";
BEGIN
	PROCESS(CLK, CLR, DISPLAY, C)
	BEGIN
		IF(CLR='1') THEN
			DISPLAY <= DIG0;
		ELSIF (CLK'EVENT AND CLK='1') THEN
			CASE C IS
				WHEN "00"=> --Retener dato
					CASE DISPLAY IS
						WHEN DIG0 => DISPLAY <= DIG0;
						WHEN DIG1 => DISPLAY <= DIG1;
						WHEN DIG2 => DISPLAY <= DIG2;
						WHEN DIG3 => DISPLAY <= DIG3;
						WHEN DIG4 => DISPLAY <= DIG4;
						WHEN DIG5 => DISPLAY <= DIG5;
						WHEN DIG6 => DISPLAY <= DIG6;
						WHEN DIG7 => DISPLAY <= DIG7;
						WHEN DIG8 => DISPLAY <= DIG8;
						WHEN DIG9 => DISPLAY <= DIG9;
						WHEN OTHERS => DISPLAY <= DIG0;
					END CASE;
				WHEN "01"=> 
					CASE DISPLAY IS
						WHEN DIG0 => DISPLAY <= DIG1;
						WHEN DIG1 => DISPLAY <= DIG2;
						WHEN DIG2 => DISPLAY <= DIG3;
						WHEN DIG3 => DISPLAY <= DIG4;
						WHEN DIG4 => DISPLAY <= DIG5;
						WHEN DIG5 => DISPLAY <= DIG6;
						WHEN DIG6 => DISPLAY <= DIG7;
						WHEN DIG7 => DISPLAY <= DIG8;
						WHEN DIG8 => DISPLAY <= DIG9;
						WHEN DIG9 => DISPLAY <= DIG0;
						WHEN OTHERS => DISPLAY <= DIG0;
					END CASE;
				WHEN "10"=> 
					CASE DISPLAY IS
						WHEN DIG0 => DISPLAY <= DIG9;
						WHEN DIG9 => DISPLAY <= DIG8;
						WHEN DIG8 => DISPLAY <= DIG7;
						WHEN DIG7 => DISPLAY <= DIG6;
						WHEN DIG6 => DISPLAY <= DIG5;
						WHEN DIG5 => DISPLAY <= DIG4;
						WHEN DIG4 => DISPLAY <= DIG3;
						WHEN DIG3 => DISPLAY <= DIG2;
						WHEN DIG2 => DISPLAY <= DIG1;
						WHEN DIG1 => DISPLAY <= DIG0;
						WHEN OTHERS => DISPLAY <= DIG0;
					END CASE;
				WHEN OTHERS => --Cargar el dato 11
					CASE E IS
						WHEN "0000" => DISPLAY <= DIG0;
						WHEN "0001" => DISPLAY <= DIG1;
						WHEN "0010" => DISPLAY <= DIG2;
						WHEN "0011" => DISPLAY <= DIG3;
						WHEN "0100" => DISPLAY <= DIG4;
						WHEN "0101" => DISPLAY <= DIG5;
						WHEN "0110" => DISPLAY <= DIG6;
						WHEN "0111" => DISPLAY <= DIG7;
						WHEN "1000" => DISPLAY <= DIG8;
						WHEN "1001" => DISPLAY <= DIG9;
						WHEN OTHERS => DISPLAY <= APAG;
					END CASE;
			END CASE;
		END IF;
	END PROCESS;
END A_CONDEC;
