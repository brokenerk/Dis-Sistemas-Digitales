module contador ( 
	clr,
	clk,
	c,
	q
	) ;

input  clr;
input  clk;
input  c;
inout [9:0] q;
