LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CONTNS IS
	PORT(CLK, CLR, C: IN STD_LOGIC;
			DISPLAY: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);

ATTRIBUTE PIN_NUMBERS OF CONTNS : ENTITY IS
"CLK:1 CLR:2 C:3 DISPLAY(0):15 DISPLAY(1):14 DISPLAY(2):22 DISPLAY(3):19 DISPLAY(4):17 DISPLAY(5):20 DISPLAY(6):18";
END ENTITY;
ARCHITECTURE A_CONTNS OF CONTNS IS
	CONSTANT H : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0001001";
	CONSTANT O : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1000000";
	CONSTANT L : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1000111";  
	CONSTANT A : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0001000";
	CONSTANT D : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100001";
	CONSTANT I : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1111001";
	CONSTANT E : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000110";
	CONSTANT Z : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100100";
BEGIN
	PROCESS(CLK, CLR, DISPLAY, C)
	BEGIN
		IF(CLR='1') THEN
			DISPLAY <= "1111111";
		ELSIF (CLK'EVENT AND CLK='1') THEN
			CASE C IS
				WHEN '0' => --HOLA
					CASE DISPLAY IS
						WHEN "1111111" => DISPLAY <= H;
						WHEN H => DISPLAY <= O;
						WHEN O => DISPLAY <= L;
						WHEN L => DISPLAY <= A;
						WHEN OTHERS => DISPLAY <= H;
					END CASE;
				WHEN OTHERS => --DIEZ
					CASE DISPLAY IS
						WHEN "1111111" => DISPLAY <= D;
						WHEN D => DISPLAY <= I;
						WHEN I => DISPLAY <= E;
						WHEN E => DISPLAY <= Z;
						WHEN OTHERS => DISPLAY <= D;
					END CASE;
			END CASE;
		END IF;
	END PROCESS;
END A_CONTNS;
