module dado ( 
	clk,
	c,
	clr,
	d
	) ;

input  clk;
input  c;
input  clr;
inout [0:6] d;
