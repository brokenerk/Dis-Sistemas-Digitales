module displays ( 
	z,
	dz
	) ;

input [1:0] z;
inout [6:0] dz;
