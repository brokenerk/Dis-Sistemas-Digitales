module ffsr ( 
	pre,
	clr,
	clk,
	s,
	r,
	q,
	nq,
	qt
	) ;

input  pre;
input  clr;
input  clk;
input  s;
input  r;
inout  q;
inout  nq;
inout  qt;
