LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG IS PORT(
	CLK, CLR, CD, CI: IN STD_LOGIC;
	C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	D: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    Q: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);

ATTRIBUTE PIN_NUMBERS OF REG: ENTITY IS
"CLK:1 C(1):2 C(0):3 D(7):4 D(6):5 D(5):6 D(4):7 D(3):8 D(2):9 D(1):10 D(0):11 Q(7):23 Q(6):22 Q(5):21 Q(4):20 Q(3):19 Q(2):18 Q(1):17 Q(0):16 CLR:15 CD:14 CI:13";


END ENTITY;
--Version 2
ARCHITECTURE A_REG OF REG IS
SIGNAL Z: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN

MUX: PROCESS(C) BEGIN
FOR I IN 7 DOWNTO 0 LOOP
	CASE C IS
		WHEN "00" => Z(I) <= Q(I);
 	    WHEN "01" => Z(I) <= D(I);
		WHEN "10" => IF (I=7) THEN
						Z(I) <= CD;
					 ELSE
					 	Z(I) <= Q(I+1);
					 END IF;
		WHEN OTHERS => IF (I=0) THEN
						Z(I) <= CI;
					 ELSE
					 	Z(I) <= Q(I-1);
					 END IF;
	END CASE;
END LOOP;
END PROCESS MUX;

REG: PROCESS (CLK, CLR) BEGIN
IF (CLR='0') THEN
	Q <= "00000000";
ELSIF (CLK'EVENT AND CLK='1') THEN
	Q <= Z;
END IF;
END PROCESS REG;
END A_REG;
