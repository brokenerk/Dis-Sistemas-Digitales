module prac1 ( 
	a,
	b,
	c,
	d,
	r,
	s,
	z,
	display
	) ;

input [1:0] a;
input [1:0] b;
input [1:0] c;
input [1:0] d;
input [1:0] r;
input [1:0] s;
inout [1:0] z;
inout [6:0] display;
