LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DISPLAYS IS PORT(
Z: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
DZ: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
);
ATTRIBUTE PIN_NUMBERS OF DISPLAYS: ENTITY IS
"Z(1):1 Z(0):2 DZ(0):20 DZ(1):19 DZ(2):18 DZ(3):17 DZ(4):16 DZ(5):15 DZ(6):14";
END ENTITY;

ARCHITECTURE A_DISPLAYS OF DISPLAYS IS 
BEGIN

DECO_Z: PROCESS (Z) BEGIN
	IF (Z="00") THEN DZ <= "0111111";
	ELSIF (Z="01") THEN DZ <= "0000110";
	ELSIF (Z="10") THEN DZ <= "1011011";
	ELSE DZ <= "1001111";
	END IF;
END PROCESS DECO_Z;
END A_DISPLAYS;
