module ffjk ( 
	pre,
	clr,
	clk,
	j,
	k,
	q,
	nq,
	qt
	) ;

input  pre;
input  clr;
input  clk;
input  j;
input  k;
inout  q;
inout  nq;
inout  qt;
