LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PRAC1 IS PORT(
A,B,C,D,R,S: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
Z: INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
DISPLAY: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
);

ATTRIBUTE PIN_NUMBERS OF PRAC1: ENTITY IS
"A(1):1 A(0):2 B(1):3 B(0):4 C(1):5 C(0):6 D(1):7 D(0):8 S(1):9 S(0):10 R(1):11 R(0):23 Z(1):22 Z(0):21 DISPLAY(2):20 DISPLAY(3):19 DISPLAY(0):18 DISPLAY(1):17 DISPLAY(4):16 DISPLAY(5):15 DISPLAY(6):14";


END ENTITY;

ARCHITECTURE A_PRAC1 OF PRAC1 IS 
SIGNAL AUX: STD_LOGIC_VECTOR (2 DOWNTO 0);

BEGIN

MUX: PROCESS (S) BEGIN
	CASE S IS
		WHEN "00" => Z <= A;
		WHEN "01" => Z <= B;
		WHEN "10" => Z <= C;
		WHEN OTHERS => Z <= D;
	END CASE;
END PROCESS MUX;

COMP: PROCESS (Z, R) BEGIN
	IF (Z=R) THEN AUX <= "100";
	ELSIF (Z>R) THEN AUX <= "010";
	ELSE AUX <= "001";
	END IF;
END PROCESS COMP;

DECO: PROCESS (AUX) BEGIN
	IF (AUX="100") THEN DISPLAY <= "1001000";
	ELSIF (AUX="010") THEN DISPLAY <= "1001100";
	ELSE DISPLAY <= "1011000";
	END IF;
END PROCESS DECO;

END A_PRAC1;
