module contreg ( 
	clk,
	clr,
	c,
	e,
	q
	) ;

input  clk;
input  clr;
input [2:0] c;
input [3:0] e;
inout [3:0] q;
