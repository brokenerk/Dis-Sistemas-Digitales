module contns ( 
	clk,
	clr,
	c,
	display
	) ;

input  clk;
input  clr;
input  c;
inout [6:0] display;
