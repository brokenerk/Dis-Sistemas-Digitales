module fft ( 
	pre,
	clr,
	clk,
	t,
	q,
	nq,
	qt
	) ;

input  pre;
input  clr;
input  clk;
input  t;
inout  q;
inout  nq;
inout  qt;
